`define TEXT 4'b1010
module test;

 initial $display("%b", `TEXT);

endmodule
